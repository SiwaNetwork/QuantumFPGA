--*****************************************************************************************
-- Project: Time Card
--
--
--
--
--
--*****************************************************************************************


--*****************************************************************************************
-- General Libraries
--*****************************************************************************************
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library TimeCardLib;
use TimeCardlib.TimeCard_Package.all;

library xil_defaultlib;
use xil_defaultlib.all;

--*****************************************************************************************
-- Entity Declaration
--*****************************************************************************************
entity TimeCardTop is
    generic (
        GoldenImage_Gen             :       boolean := false
    );
    port (
        -- System 
        Mhz10ClkDcxo1_ClkIn         : in    std_logic;
            
        RstN_RstIn                  : in    std_logic;
        
        -- MAC RF Out Clock
        Mhz10Clk0_ClkIn             : in    std_logic;
        Mhz10Clk1_ClkIn             : in    std_logic;
        
        --GTP Clock
        Mhz125ClkP_ClkIn            : in    std_logic;
        Mhz125ClkN_ClkIn            : in    std_logic;
        
        --200MHz Clock
        Mhz200ClkP_ClkIn            : in    std_logic;
        Mhz200ClkN_ClkIn            : in    std_logic; 
        
        Led_DatOut                  : out   std_logic_vector(3 downto 0);
        Key_DatIn                   : in    std_logic_vector(1 downto 0);
   
        EepromWp_DatOut             : out   std_logic;
   
        -----------------------------------------------------------------
        -- QSPI Flash Inputs/Outputs
        -----------------------------------------------------------------
        SpiFlashDq0_DatInOut        : inout std_logic;
        SpiFlashDq1_DatInOut        : inout std_logic;
        SpiFlashDq2_DatInOut        : inout std_logic;
        SpiFlashDq3_DatInOut        : inout std_logic;
        SpiFlashCsN_EnaOut          : out   std_logic;
        
        -----------------------------------------------------------------
        -- SMA Inputs/Outputs
        -----------------------------------------------------------------
        SmaIn1_DatIn                : in    std_logic;      -- ANT1
        SmaIn2_DatIn                : in    std_logic;      -- ANT2
        SmaIn3_DatIn                : in    std_logic;      -- ANT3
        SmaIn4_DatIn                : in    std_logic;      -- ANT4
        
        SmaOut1_DatOut              : out   std_logic;      -- ANT1
        SmaOut2_DatOut              : out   std_logic;      -- ANT2
        SmaOut3_DatOut              : out   std_logic;      -- ANT3
        SmaOut4_DatOut              : out   std_logic;      -- ANT4
        
        Sma1InBufEnableN_EnOut      : out   std_logic;
        Sma2InBufEnableN_EnOut      : out   std_logic;
        Sma3InBufEnableN_EnOut      : out   std_logic;
        Sma4InBufEnableN_EnOut      : out   std_logic;
        
        Sma1OutBufEnableN_EnOut     : out   std_logic;
        Sma2OutBufEnableN_EnOut     : out   std_logic;
        Sma3OutBufEnableN_EnOut     : out   std_logic;
        Sma4OutBufEnableN_EnOut     : out   std_logic;
        
        -----------------------------------------------------------------
        -- I2C
        -----------------------------------------------------------------
        I2cScl_ClkInOut             : inout std_logic;
        I2cSda_DatInOut             : inout std_logic;
        
        -----------------------------------------------------------------
        -- UART1
        -----------------------------------------------------------------
        Uart1TxDat_DatOut           : out   std_logic;
        Uart1RxDat_DatIn            : in    std_logic;
        
        -----------------------------------------------------------------
        -- GNSS
        -----------------------------------------------------------------
        UartGnss1TxDat_DatOut       : out   std_logic;
        UartGnss1RxDat_DatIn        : in    std_logic;
        Gnss1Tp_DatIn               : in    std_logic_vector(1 downto 0);
        Gnss1RstN_RstOut            : out   std_logic;
        
        UartGnss2TxDat_DatOut       : out   std_logic;
        UartGnss2RxDat_DatIn        : in    std_logic;
        Gnss2Tp_DatIn               : in    std_logic_vector(1 downto 0);
        Gnss2RstN_RstOut            : out   std_logic;
        
        -----------------------------------------------------------------
        --MAC
        -----------------------------------------------------------------
        MacTxDat_DatInOut           : inout std_logic;
        MacRxDat_DatInOut           : inout std_logic;
        
        MacFreqControl_DatOut       : out   std_logic;
        MacAlarm_DatIn              : in    std_logic;
        MacBite_DatIn               : in    std_logic;
        
        MacUsbPower_EnOut           : out   std_logic;
        MacUsbP_DatOut              : out   std_logic;
        MacUsbN_DatOut              : out   std_logic;
        
        MacPps_EvtIn                : in    std_logic;
        MacPps0_EvtOut              : out   std_logic;
        MacPps1_EvtOut              : out   std_logic;

        -----------------------------------------------------------------
        --PCIe
        -----------------------------------------------------------------
        PciePerst_RstIn             : in    std_logic;
        PcieRefClkP_ClkIn           : in    std_logic;
        PcieRefClkN_ClkIn           : in    std_logic;
        pcie_7x_mgt_0_rxn           : in    std_logic_vector(0 downto 0);
        pcie_7x_mgt_0_rxp           : in    std_logic_vector(0 downto 0);
        pcie_7x_mgt_0_txn           : out   std_logic_vector(0 downto 0);
        pcie_7x_mgt_0_txp           : out   std_logic_vector(0 downto 0)
    );
end TimeCardTop;

--*****************************************************************************************
-- Architecture Declaration
--*****************************************************************************************
architecture TimeCardTop_Arch of TimeCardTop is
    --*************************************************************************************
    -- Component Definitions
    --*************************************************************************************
    component Bufio
        port (
            i                           : in    std_logic; 
            o                           : out   std_logic
        );
    end component Bufio;    
    
    
    component Bufg
        port (
            i                           : in    std_logic; 
            o                           : out   std_logic
        );
    end component Bufg;    
        
    component Bufr is
        port (
            o                           : out std_logic;
            ce                          : in std_logic;
            clr                         : in std_logic;
            i                           : in std_logic
        );
    end component Bufr;
    
    component Ibufds is
        port (
            i                           : in    std_logic;
            ib                          : in    std_logic;
            o                           : out   std_logic
        );
    end component Ibufds;
    
    component Obufds is
        port (
            o                           : out   std_logic;
            ob                          : out   std_logic;
            i                           : in    std_logic
        );
    end component Obufds;

    component litepcie_core is
    port (
        clk                         	: out 	std_logic;
        rst                         	: out 	std_logic;
			
        ptm_time_clk                	: in	std_logic;
        ptm_time_rst                	: in	std_logic;
        ptm_time_ns                 	: in	std_logic_vector(63 downto 0);
			
        pcie_rst_n                  	: in	std_logic;
        pcie_clk_p                  	: in	std_logic;
        pcie_clk_n                  	: in	std_logic;
        pcie_rx_p                   	: in	std_logic;
        pcie_rx_n                   	: in	std_logic;
        pcie_tx_p                   	: out 	std_logic;
        pcie_tx_n                   	: out 	std_logic;
						
        mmap_axi_lite_awvalid       	: out 	std_logic;
        mmap_axi_lite_awready       	: in 	std_logic;
        mmap_axi_lite_awaddr        	: out 	std_logic_vector(31 downto 0);
        mmap_axi_lite_awprot        	: out 	std_logic_vector(2 downto 0);
        mmap_axi_lite_wvalid        	: out 	std_logic;
        mmap_axi_lite_wready        	: in 	std_logic;
        mmap_axi_lite_wdata         	: out 	std_logic_vector(31 downto 0);
        mmap_axi_lite_wstrb         	: out 	std_logic_vector(3 downto 0);
        mmap_axi_lite_bvalid        	: in 	std_logic;
        mmap_axi_lite_bready        	: out 	std_logic;
        mmap_axi_lite_bresp         	: in 	std_logic_vector(1 downto 0);
        mmap_axi_lite_arvalid       	: out 	std_logic;
        mmap_axi_lite_arready       	: in 	std_logic;
        mmap_axi_lite_araddr        	: out 	std_logic_vector(31 downto 0);
        mmap_axi_lite_arprot        	: out 	std_logic_vector(2 downto 0);
        mmap_axi_lite_rvalid        	: in 	std_logic;
        mmap_axi_lite_rready        	: out 	std_logic;
        mmap_axi_lite_rresp         	: in 	std_logic_vector(1 downto 0);
        mmap_axi_lite_rdata         	: in 	std_logic_vector(31 downto 0);
        mmap_slave_axi_lite_awvalid		: in	std_logic;
        mmap_slave_axi_lite_awready		: out 	std_logic;
        mmap_slave_axi_lite_awaddr 		: in	std_logic_vector(31 downto 0);
        mmap_slave_axi_lite_awprot 		: in	std_logic_vector(2 downto 0);
        mmap_slave_axi_lite_wvalid 		: in	std_logic;
        mmap_slave_axi_lite_wready 		: out 	std_logic;
        mmap_slave_axi_lite_wdata  		: in	std_logic_vector(31 downto 0);
        mmap_slave_axi_lite_wstrb  		: in	std_logic_vector(3 downto 0);
        mmap_slave_axi_lite_bvalid 		: out 	std_logic;
        mmap_slave_axi_lite_bready 		: in	std_logic;
        mmap_slave_axi_lite_bresp  		: out 	std_logic_vector(1 downto 0);
        mmap_slave_axi_lite_arvalid		: in	std_logic;
        mmap_slave_axi_lite_arready		: out 	std_logic;
        mmap_slave_axi_lite_araddr 		: in	std_logic_vector(31 downto 0);
        mmap_slave_axi_lite_arprot 		: in	std_logic_vector(2 downto 0);
        mmap_slave_axi_lite_rvalid 		: out 	std_logic;
        mmap_slave_axi_lite_rready 		: in	std_logic;
        mmap_slave_axi_lite_rresp  		: out 	std_logic_vector(1 downto 0);
        mmap_slave_axi_lite_rdata  		: out 	std_logic_vector(31 downto 0);
		
        msi_irqs                    	: in	std_logic_vector(31 downto 0 )
    );
    end component litepcie_core;

    
    --*************************************************************************************
    -- Procedure Definitions
    --*************************************************************************************

    --*************************************************************************************
    -- Function Definitions
    --*************************************************************************************

    --*************************************************************************************
    -- Constant Definitions
    --*************************************************************************************
    constant ClkPeriodNanosecond_Con    : natural := 20;
	
    --*************************************************************************************
    -- Type Definitions
    --*************************************************************************************

    --*************************************************************************************
    -- Signal Definitions
    --*************************************************************************************
    
    -- Rst & Clk
    signal PciePerstN_Rst               : std_logic;
    
    signal Mhz10Clk0_Clk                : std_logic;
 
    signal Mhz10ClkDcxo1_Clk            : std_logic;
    signal Mhz10ClkDcxo2_Clk            : std_logic;
    
    signal Mhz50Clk_Clk                 : std_logic;
    signal Mhz50RstN_Rst                : std_logic;
    
    signal Mhz50Clk_Clk_0               : std_logic;
    signal Mhz50RstN_Rst_0              : std_logic;
    
    signal Mhz62_5Clk_Clk               : std_logic;
    signal Mhz62_5Rst_Rst               : std_logic;
    signal Mhz62_5RstN_Rst              : std_logic;
    
    signal RstCount_CntReg              : natural := 0;
    
    -- Led
    signal BlinkingLed_DatReg           : std_logic;
    signal BlinkingLedCount_CntReg      : natural;
    
    signal BlinkingLed2_DatReg          : std_logic;
    signal BlinkingLed2Count_CntReg     : natural;
    
    -- Time 
    signal time_out_clock_nanosecond    : std_logic_vector(31 downto 0);
    signal time_out_clock_second        : std_logic_vector(31 downto 0);
    signal time_out_clock_timejump      : std_logic;
    signal time_out_clock_valid         : std_logic;
    
    signal ptm_time_clk                 : std_logic;
    signal ptm_time_rst                 : std_logic;
    signal ptm_time_ns                  : std_logic_vector(63 downto 0);
    
    signal GnssDataOe_EnaReg            : std_logic;
    
    signal Ext_DatIn                    : std_logic_vector(1 downto 0);
    signal Ext_DatOut                   : std_logic_vector(6 downto 0);
    
    signal Pps_EvtOut                   : std_logic;

    signal MacPps0_Evt                  : std_logic;
    signal MacPps1_Evt                  : std_logic;
    signal GpioGnss_DatOut              : std_logic_vector(1 downto 0);
    
    signal UartGnss1TxDat_Dat           : std_logic;
    signal UartGnss2TxDat_Dat           : std_logic;
        
    signal StartUpIo_cfgclk             : std_logic;
    signal StartUpIo_cfgmclk            : std_logic;
    signal StartUpIo_preq               : std_logic;
    
    -- SMA Connector / Buffers
    signal SmaIn1_En                    : std_logic;
    signal SmaIn2_En                    : std_logic;
    signal SmaIn3_En                    : std_logic;
    signal SmaIn4_En                    : std_logic;
        
    signal SmaOut1_En                   : std_logic;
    signal SmaOut2_En                   : std_logic;
    signal SmaOut3_En                   : std_logic;
    signal SmaOut4_En                   : std_logic;
    
    signal SpiFlashCsN_Ena              : std_logic;
    
    signal GoldenImageN_Ena             : std_logic;
    
    signal Clk_RxSda_i                  : std_logic;
    signal Clk_RxSda_o                  : std_logic;
    signal Clk_RxSda_t                  : std_logic;
    signal Clk_TxScl_i                  : std_logic;
    signal Clk_TxScl_o                  : std_logic;
    signal Clk_TxScl_t                  : std_logic;
    
    signal Msi_Dat                      : std_logic_vector(31 downto 0) := (others => '0');

    -- AXI  
    signal mmap_axi_lite_awvalid        : std_logic_vector(0 downto 0);
    signal awvalid                      : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_awready        : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_awaddr         : std_logic_vector(31 downto 0);
    signal awaddr                       : std_logic_vector(31 downto 0);
    signal mmap_axi_lite_awprot         : std_logic_vector(2 downto 0);
    signal mmap_axi_lite_wvalid         : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_wready         : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_wdata          : std_logic_vector(31 downto 0);
    signal mmap_axi_lite_wstrb          : std_logic_vector(3 downto 0);
    signal mmap_axi_lite_bvalid         : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_bready         : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_bresp          : std_logic_vector(1 downto 0);
    signal mmap_axi_lite_arvalid        : std_logic_vector(0 downto 0);
    signal arvalid                      : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_arready        : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_araddr         : std_logic_vector(31 downto 0);
    signal araddr                       : std_logic_vector(31 downto 0);
    signal mmap_axi_lite_arprot         : std_logic_vector(2 downto 0);
    signal mmap_axi_lite_rvalid         : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_rready         : std_logic_vector(0 downto 0);
    signal mmap_axi_lite_rresp          : std_logic_vector(1 downto 0);
    signal mmap_axi_lite_rdata          : std_logic_vector(31 downto 0);
    
    signal mmap_slave_axi_lite_awvalid  : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_awready  : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_awaddr   : std_logic_vector(31 downto 0);
    signal mmap_slave_axi_lite_awprot   : std_logic_vector(2 downto 0);
    signal mmap_slave_axi_lite_wvalid   : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_wready   : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_wdata    : std_logic_vector(31 downto 0);
    signal mmap_slave_axi_lite_wstrb    : std_logic_vector(3 downto 0);
    signal mmap_slave_axi_lite_bvalid   : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_bready   : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_bresp    : std_logic_vector(1 downto 0);
    signal mmap_slave_axi_lite_arvalid  : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_arready  : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_araddr   : std_logic_vector(31 downto 0);
    signal mmap_slave_axi_lite_arprot   : std_logic_vector(2 downto 0);
    signal mmap_slave_axi_lite_rvalid   : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_rready   : std_logic_vector(0 downto 0);
    signal mmap_slave_axi_lite_rresp    : std_logic_vector(1 downto 0);
    signal mmap_slave_axi_lite_rdata    : std_logic_vector(31 downto 0);
    
--*****************************************************************************************
-- Architecture Implementation
--*****************************************************************************************
begin
    --*************************************************************************************
    -- Concurrent Statements
    --*************************************************************************************
    
    -- CLK UART and CLK I2C share the same pins (it is configurable which interface is active)
    Clk_RxSda_i <= MacRxDat_DatInOut;
    MacRxDat_DatInOut <= Clk_RxSda_o when (Clk_RxSda_t = '0') else 'Z';
    
    Clk_TxScl_i <= MacTxDat_DatInOut;
    MacTxDat_DatInOut <= Clk_TxScl_o when (Clk_TxScl_t = '0') else 'Z';
    
    -- SMA
    Sma1InBufEnableN_EnOut <= not SmaIn1_En;
    Sma2InBufEnableN_EnOut <= not SmaIn2_En;
    Sma3InBufEnableN_EnOut <= not SmaIn3_En;
    Sma4InBufEnableN_EnOut <= not SmaIn4_En;
    
    Sma1OutBufEnableN_EnOut <= not SmaOut1_En;
    Sma2OutBufEnableN_EnOut <= not SmaOut2_En;
    Sma3OutBufEnableN_EnOut <= not SmaOut3_En;
    Sma4OutBufEnableN_EnOut <= not SmaOut4_En;
    
    
    GoldenImageN_Ena <= '0' when GoldenImage_Gen = true else '1';
    
    PciePerstN_Rst <= PciePerst_RstIn;
    
    Ext_DatIn <= Key_DatIn;
    
    Led_DatOut(3) <= MacPps_EvtIn;          -- Ext_DatOut(3);
    Led_DatOut(2) <= Pps_EvtOut;            -- Ext_DatOut(2);
    Led_DatOut(1) <= BlinkingLed2_DatReg;   -- Ext_DatOut(1);
    Led_DatOut(0) <= BlinkingLed_DatReg;    -- Ext_DatOut(0);
    
    EepromWp_DatOut <= Ext_DatOut(4);
    
    -- GNSS Outputs
    Gnss1RstN_RstOut <= not GpioGnss_DatOut(0);
    Gnss2RstN_RstOut <= not GpioGnss_DatOut(1);
    
    -- Wait 1s until enable Gnss Uart Tx Output
    UartGnss1TxDat_DatOut <= 'Z' when GnssDataOe_EnaReg = '0' else UartGnss1TxDat_Dat;
    UartGnss2TxDat_DatOut <= 'Z' when GnssDataOe_EnaReg = '0' else UartGnss2TxDat_Dat;
    
    -- SPI Flash
    SpiFlashCsN_EnaOut <= SpiFlashCsN_Ena;
    
    -- MAC
    MacFreqControl_DatOut <= '0';
    MacUsbPower_EnOut <= '0';
    
    --! unused uart
    Uart1TxDat_DatOut <= '0'; --! unused

    --*************************************************************************************
    -- Procedural Statements
    --*************************************************************************************
    BlinkingLed_Prc : process(Mhz50RstN_Rst, Mhz50Clk_Clk) is
    begin
        if (Mhz50RstN_Rst = '0') then
            BlinkingLed_DatReg <= '0';
            BlinkingLedCount_CntReg <= 0;
        elsif ((Mhz50Clk_Clk'event) and (Mhz50Clk_Clk = '1')) then
            if (BlinkingLedCount_CntReg < 250000000) then
                BlinkingLedCount_CntReg <= BlinkingLedCount_CntReg + ClkPeriodNanosecond_Con;
            else
                BlinkingLed_DatReg <= (not BlinkingLed_DatReg);
                BlinkingLedCount_CntReg <= 0;
            end if;
        end if;
    end process BlinkingLed_Prc;
    
    BlinkingLed2_Prc : process(Mhz62_5RstN_Rst, Mhz62_5Clk_Clk) is
    begin
        if (Mhz62_5RstN_Rst = '0') then
            BlinkingLed2_DatReg <= '0';
            BlinkingLed2Count_CntReg <= 0;
        elsif ((Mhz62_5Clk_Clk'event) and (Mhz62_5Clk_Clk = '1')) then
            if (BlinkingLed2Count_CntReg < 200000000) then
                BlinkingLed2Count_CntReg <= BlinkingLed2Count_CntReg + ClkPeriodNanosecond_Con;
            else
                BlinkingLed2_DatReg <= (not BlinkingLed2_DatReg);
                BlinkingLed2Count_CntReg <= 0;
            end if;
        end if;
    end process BlinkingLed2_Prc;
    
    Rst_Prc : process(Mhz50RstN_Rst, Mhz50Clk_Clk) is
    begin
        if (Mhz50RstN_Rst = '0') then
            GnssDataOe_EnaReg <= '0';
            RstCount_CntReg <= 0;
        elsif ((Mhz50Clk_Clk'event) and (Mhz50Clk_Clk = '1')) then
            if (RstCount_CntReg < 2000000000) then
                RstCount_CntReg <= RstCount_CntReg + ClkPeriodNanosecond_Con;
                if (RstCount_CntReg < 1000000000) then -- 1000ms
                    GnssDataOe_EnaReg <= '0';
                else
                    GnssDataOe_EnaReg <= '1';
                end if;
            else
                RstCount_CntReg <= RstCount_CntReg;
                GnssDataOe_EnaReg <= '1';
            end if;
        end if;
    end process Rst_Prc;
    
    --*************************************************************************************
    -- Instantiation and Port mapping
    --*************************************************************************************
    
    MacPps0_EvtOut <= MacPps0_Evt;
    MacPps1_EvtOut <= MacPps1_Evt;
    
    -- MacUsb_Inst: component Obufds 
    -- port map(
        -- o                           => MacUsbP_DatOut,
        -- ob                          => MacUsbN_DatOut,
        -- i                           => '0'
    -- );
    MacUsbP_DatOut <= '0';
    MacUsbN_DatOut <= '0';
       
    
    BufrClk0_Inst : Bufr   
    port map (  
        ce                              => '1',
        clr                             => '0',
        i                               => Mhz10Clk0_ClkIn,
        o                               => Mhz10Clk0_Clk
    );  
    
    BufrDcxo1_Inst : Bufr   
    port map (
        ce                              => '1',
        clr                             => '0',
        i                               => Mhz10ClkDcxo1_ClkIn,
        o                               => Mhz10ClkDcxo1_Clk
    );   
   
    -- BufrDcxo2_Inst : Bufr   
    -- port map (
        -- ce                              => '1',
        -- clr                             => '0',
        -- i                               => Mhz10ClkDcxo2_ClkIn,
        -- o                               => Mhz10ClkDcxo2_Clk
    -- );      

    Mhz62_5RstN_Rst <= not Mhz62_5Rst_Rst;

    ptm_time_clk <= Mhz50Clk_Clk;
    ptm_time_rst <= not Mhz50RstN_Rst;
    ptm_time_ns <= std_logic_vector(resize(unsigned(time_out_clock_second(31 downto 0)) * to_unsigned(SecondNanoseconds_Con, 32) + unsigned(time_out_clock_nanosecond), 64));

    PciE: litepcie_core
    port map (
        clk                             => Mhz62_5Clk_Clk,
        rst                             => Mhz62_5Rst_Rst,
        pcie_rst_n                      => PciePerstN_Rst,
        
        ptm_time_clk                    => ptm_time_clk,
        ptm_time_rst                    => ptm_time_rst,
        ptm_time_ns                     => ptm_time_ns,
        
        -- pcie_rst_n                      => '0',
        pcie_clk_p                      => PcieRefClkP_ClkIn,
        pcie_clk_n                      => PcieRefClkN_ClkIn,
        pcie_rx_p                       => pcie_7x_mgt_0_rxp(0),
        pcie_rx_n                       => pcie_7x_mgt_0_rxn(0),
        pcie_tx_p                       => pcie_7x_mgt_0_txp(0),
        pcie_tx_n                       => pcie_7x_mgt_0_txn(0),
                
        mmap_axi_lite_awvalid           => mmap_axi_lite_awvalid(0),  
        mmap_axi_lite_awready           => mmap_axi_lite_awready(0),  
        mmap_axi_lite_awaddr            => mmap_axi_lite_awaddr,      
        mmap_axi_lite_awprot            => mmap_axi_lite_awprot,      
        mmap_axi_lite_wvalid            => mmap_axi_lite_wvalid(0),   
        mmap_axi_lite_wready            => mmap_axi_lite_wready(0),   
        mmap_axi_lite_wdata             => mmap_axi_lite_wdata,       
        mmap_axi_lite_wstrb             => mmap_axi_lite_wstrb,       
        mmap_axi_lite_bvalid            => mmap_axi_lite_bvalid(0),   
        mmap_axi_lite_bready            => mmap_axi_lite_bready(0),   
        mmap_axi_lite_bresp             => mmap_axi_lite_bresp,       
        mmap_axi_lite_arvalid           => mmap_axi_lite_arvalid(0),  
        mmap_axi_lite_arready           => mmap_axi_lite_arready(0),  
        mmap_axi_lite_araddr            => mmap_axi_lite_araddr,      
        mmap_axi_lite_arprot            => mmap_axi_lite_arprot,      
        mmap_axi_lite_rvalid            => mmap_axi_lite_rvalid(0),   
        mmap_axi_lite_rready            => mmap_axi_lite_rready(0),   
        mmap_axi_lite_rresp             => mmap_axi_lite_rresp,       
        mmap_axi_lite_rdata             => mmap_axi_lite_rdata,       
    
        mmap_slave_axi_lite_awvalid     => mmap_slave_axi_lite_awvalid(0),  
        mmap_slave_axi_lite_awready     => mmap_slave_axi_lite_awready(0),  
        mmap_slave_axi_lite_awaddr      => mmap_slave_axi_lite_awaddr,      
        mmap_slave_axi_lite_awprot      => mmap_slave_axi_lite_awprot,      
        mmap_slave_axi_lite_wvalid      => mmap_slave_axi_lite_wvalid(0),   
        mmap_slave_axi_lite_wready      => mmap_slave_axi_lite_wready(0),   
        mmap_slave_axi_lite_wdata       => mmap_slave_axi_lite_wdata,       
        mmap_slave_axi_lite_wstrb       => mmap_slave_axi_lite_wstrb,       
        mmap_slave_axi_lite_bvalid      => mmap_slave_axi_lite_bvalid(0),   
        mmap_slave_axi_lite_bready      => mmap_slave_axi_lite_bready(0),   
        mmap_slave_axi_lite_bresp       => mmap_slave_axi_lite_bresp,       
        mmap_slave_axi_lite_arvalid     => mmap_slave_axi_lite_arvalid(0),  
        mmap_slave_axi_lite_arready     => mmap_slave_axi_lite_arready(0),  
        mmap_slave_axi_lite_araddr      => mmap_slave_axi_lite_araddr,      
        mmap_slave_axi_lite_arprot      => mmap_slave_axi_lite_arprot,      
        mmap_slave_axi_lite_rvalid      => mmap_slave_axi_lite_rvalid(0),   
        mmap_slave_axi_lite_rready      => mmap_slave_axi_lite_rready(0),   
        mmap_slave_axi_lite_rresp       => mmap_slave_axi_lite_rresp,       
        mmap_slave_axi_lite_rdata       => mmap_slave_axi_lite_rdata,       

        msi_irqs                        => Msi_Dat
    );
    
    Bd_Inst : entity xil_defaultlib.TimeCard_wrapper
    port map (
        Mhz200Clk_ClkIn_clk_n       => Mhz200ClkN_ClkIn,
        Mhz200Clk_ClkIn_clk_p       => Mhz200ClkP_ClkIn,
        
        Mhz10ClkMac_ClkIn           => Mhz10Clk0_Clk,
        Mhz10ClkSma_ClkIn           => SmaIn1_DatIn,
        Mhz10ClkDcxo1_ClkIn         => Mhz10ClkDcxo1_Clk,
        Mhz10ClkDcxo2_ClkIn         => '0',
        
        ResetN_RstIn                => RstN_RstIn,
        GoldenImageN_EnaIn          => GoldenImageN_Ena,
       
        -- Internal 50MHz (does no change on clock source switch)
        Mhz50Clk_ClkOut_0           => Mhz50Clk_Clk_0,
        Reset50MhzN_RstOut_0(0)     => Mhz50RstN_Rst_0,    
        
        Mhz50Clk_ClkOut             => Mhz50Clk_Clk,
        Reset50MhzN_RstOut(0)       => Mhz50RstN_Rst,       

--!        Mhz62_5Clk_ClkOut           => Mhz62_5Clk_Clk,
--!        Reset62_5MhzN_RstOut(0)     => Mhz62_5RstN_Rst,

        InHoldover_DatOut           => open,
        InSync_DatOut               => open,
        
        Ext_DatIn_tri_i             => Ext_DatIn,
        Ext_DatOut                  => Ext_DatOut,
        
        I2c_scl_io                  => I2cScl_ClkInOut,
        I2c_sda_io                  => I2cSda_DatInOut,
        
        SpiFlash_io0_io             => SpiFlashDq0_DatInOut,
        SpiFlash_io1_io             => SpiFlashDq1_DatInOut,
        SpiFlash_io2_io             => SpiFlashDq2_DatInOut,
        SpiFlash_io3_io             => SpiFlashDq3_DatInOut,
        SpiFlash_ss_io(0)           => SpiFlashCsN_Ena,
        
        StartUpIo_cfgclk            => StartUpIo_cfgclk,
        StartUpIo_cfgmclk           => StartUpIo_cfgmclk,
        StartUpIo_preq              => StartUpIo_preq,
        
        GpioGnss_DatOut_tri_o       => GpioGnss_DatOut,

        GpioMac_DatIn_tri_i(0)      => MacAlarm_DatIn,
        GpioMac_DatIn_tri_i(1)      => MacBite_DatIn,
        
        SmaIn1_DatIn                => SmaIn1_DatIn,
        SmaIn1_EnOut                => SmaIn1_En,
        SmaIn2_DatIn                => SmaIn2_DatIn,
        SmaIn2_EnOut                => SmaIn2_En,
        SmaIn3_DatIn                => SmaIn3_DatIn,
        SmaIn3_EnOut                => SmaIn3_En,
        SmaIn4_DatIn                => SmaIn4_DatIn,
        SmaIn4_EnOut                => SmaIn4_En,
        
        SmaOut1_DatOut              => SmaOut1_DatOut,
        SmaOut1_EnOut               => SmaOut1_En,
        SmaOut2_DatOut              => SmaOut2_DatOut,
        SmaOut2_EnOut               => SmaOut2_En,
        SmaOut3_DatOut              => SmaOut3_DatOut,
        SmaOut3_EnOut               => SmaOut3_En,
        SmaOut4_DatOut              => SmaOut4_DatOut,
        SmaOut4_EnOut               => SmaOut4_En,

        PpsGnss1_EvtIn              => Gnss1Tp_DatIn(0),
        PpsGnss2_EvtIn              => Gnss2Tp_DatIn(0),
        Pps_EvtOut                  => Pps_EvtOut,
        
        MacPps_EvtIn                => MacPps_EvtIn,
        MacPps0_EvtOut              => MacPps0_Evt,
        MacPps1_EvtOut              => MacPps1_Evt,

        UartGnss1Rx_DatIn           => UartGnss1RxDat_DatIn,
        UartGnss1Tx_DatOut          => UartGnss1TxDat_Dat,
        
        UartGnss2Rx_DatIn           => UartGnss2RxDat_DatIn,
        UartGnss2Tx_DatOut          => UartGnss2TxDat_Dat,
        
        time_out_nanosecond         => time_out_clock_nanosecond,
        time_out_second             => time_out_clock_second,
        time_out_timejump           => time_out_clock_timejump,
        time_out_valid              => time_out_clock_valid,
        
        Clk_RxSda_DatIn             => Clk_RxSda_i,
        Clk_RxSda_DatOut            => Clk_RxSda_o,
        Clk_RxSdaT_EnaOut           => Clk_RxSda_t,
        Clk_TxSclT_EnaOut           => Clk_TxScl_t,
        Clk_TxScl_DatIn             => Clk_TxScl_i,
        Clk_TxScl_DatOut            => Clk_TxScl_o,

        Mhz62_5Clk_ClkIn            => Mhz62_5Clk_Clk,
        PciePerstN_RstIn            => PciePerstN_Rst,

        -- PCIe MMAP 
        mmap_axi_lite_awaddr         => awaddr,
        -- mmap_axi_lite_awaddr         => mmap_axi_lite_awaddr,
        mmap_axi_lite_awprot         => mmap_axi_lite_awprot,
        mmap_axi_lite_awvalid        => awvalid,
        mmap_axi_lite_awready        => mmap_axi_lite_awready,
        mmap_axi_lite_wdata          => mmap_axi_lite_wdata,
        mmap_axi_lite_wstrb          => mmap_axi_lite_wstrb,
        mmap_axi_lite_wvalid         => mmap_axi_lite_wvalid,
        mmap_axi_lite_wready         => mmap_axi_lite_wready,
        mmap_axi_lite_bresp          => mmap_axi_lite_bresp,
        mmap_axi_lite_bvalid         => mmap_axi_lite_bvalid,
        mmap_axi_lite_bready         => mmap_axi_lite_bready,
        mmap_axi_lite_araddr         => araddr,
        -- mmap_axi_lite_araddr         => mmap_axi_lite_araddr,
        mmap_axi_lite_arprot         => mmap_axi_lite_arprot,
        mmap_axi_lite_arvalid        => arvalid,
        mmap_axi_lite_arready        => mmap_axi_lite_arready,
        mmap_axi_lite_rdata          => mmap_axi_lite_rdata,
        mmap_axi_lite_rresp          => mmap_axi_lite_rresp,
        mmap_axi_lite_rvalid         => mmap_axi_lite_rvalid,
        mmap_axi_lite_rready         => mmap_axi_lite_rready,
        
        -- Interrupts to PCIe
        Msi_DatOut                  => Msi_Dat(19 downto 0),
        -- PCIe slave
        M_Pcie_Ctl_awaddr           => mmap_slave_axi_lite_awaddr,
        M_Pcie_Ctl_awprot           => mmap_slave_axi_lite_awprot,
        M_Pcie_Ctl_awvalid          => mmap_slave_axi_lite_awvalid,
        M_Pcie_Ctl_awready          => mmap_slave_axi_lite_awready,
        M_Pcie_Ctl_wdata            => mmap_slave_axi_lite_wdata,
        M_Pcie_Ctl_wstrb            => mmap_slave_axi_lite_wstrb,
        M_Pcie_Ctl_wvalid           => mmap_slave_axi_lite_wvalid,
        M_Pcie_Ctl_wready           => mmap_slave_axi_lite_wready,
        M_Pcie_Ctl_bresp            => mmap_slave_axi_lite_bresp,
        M_Pcie_Ctl_bvalid           => mmap_slave_axi_lite_bvalid,
        M_Pcie_Ctl_bready           => mmap_slave_axi_lite_bready,
        M_Pcie_Ctl_araddr           => mmap_slave_axi_lite_araddr,
        M_Pcie_Ctl_arprot           => mmap_slave_axi_lite_arprot,
        M_Pcie_Ctl_arvalid          => mmap_slave_axi_lite_arvalid,
        M_Pcie_Ctl_arready          => mmap_slave_axi_lite_arready,
        M_Pcie_Ctl_rdata            => mmap_slave_axi_lite_rdata,
        M_Pcie_Ctl_rresp            => mmap_slave_axi_lite_rresp,
        M_Pcie_Ctl_rvalid           => mmap_slave_axi_lite_rvalid,
        M_Pcie_Ctl_rready           => mmap_slave_axi_lite_rready
    );

    awaddr <= "0000000" & mmap_axi_lite_awaddr(24 downto 0);
    araddr <= "0000000" & mmap_axi_lite_araddr(24 downto 0);
    
    awvalid(0) <= mmap_axi_lite_awvalid(0) and mmap_axi_lite_awaddr(25);
    arvalid(0) <= mmap_axi_lite_arvalid(0) and mmap_axi_lite_araddr(25);
    
end TimeCardTop_Arch;
