--*****************************************************************************************
-- Проект: Time Card
--
--
--
--
--
--*****************************************************************************************

--*****************************************************************************************
-- Общие библиотеки
--*****************************************************************************************
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

--*****************************************************************************************
-- Специфические библиотеки
--*****************************************************************************************

--*****************************************************************************************
-- Объявление сущности
--*****************************************************************************************
entity SinglePulseIrq is

    port (
        -- System
        SysClk_ClkIn                    : in    std_logic;
        SysRstN_RstIn                   : in    std_logic;

        -- Interrupt input         
        IrqIn_DatIn                     : in    std_logic;

        -- Interrupt output         
        IrqOut_DatOut                   : out   std_logic
    );
end entity SinglePulseIrq;


--*****************************************************************************************
-- Объявление архитектуры
--*****************************************************************************************
architecture SinglePulseIrq_Arch of SinglePulseIrq is
    --*************************************************************************************
    -- Определения процедур
    --*************************************************************************************

    --*************************************************************************************
    -- Определения функций
    --*************************************************************************************

    --*************************************************************************************
    -- Определения констант
    --*************************************************************************************

    --*************************************************************************************
    -- Определения типов
    --*************************************************************************************

    --*************************************************************************************
    -- Определения сигналов
    --*************************************************************************************
    signal IrqIn_DatReg                     : std_logic;
    signal IrqIn_DatOutReg                  : std_logic;
    
    --*****************************************************************************************
-- Реализация архитектуры
--*****************************************************************************************
begin

    --*************************************************************************************
    -- Конкурентные операторы
    --*************************************************************************************
    IrqOut_DatOut <= IrqIn_DatOutReg;
    
    --*************************************************************************************
    -- Процедурные операторы
    --*************************************************************************************
    SignlePulsIrq_Prc : process(SysClk_ClkIn, SysRstN_RstIn) is
    begin
        if (SysRstN_RstIn = '0') then
            IrqIn_DatReg <= '0';
            IrqIn_DatOutReg <= '0';
        elsif ((SysClk_ClkIn'event) and (SysClk_ClkIn = '1')) then
            IrqIn_DatReg <= IrqIn_DatIn;
            IrqIn_DatOutReg <= '0';
     
            if (IrqIn_DatIn = '1' and IrqIn_DatReg = '0') then
                IrqIn_DatOutReg <= '1';
            end if;
        end if;
    end process SignlePulsIrq_Prc;
    
    --*************************************************************************************
    -- Инстанцирование и отображение портов
    --*************************************************************************************
        
end architecture SinglePulseIrq_Arch;